localparam period = 1.43;
localparam halfperiod = period/2;
parameter width1 = 8;
parameter width2 = 8;
parameter outwidth = 16;
